// $Id: $
// File name:   rcv_block.sv
// Created:     2/11/2016
// Author:      Chongjin Chua
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: rcv_block.sv

module rcv_block
  (
   input wire clk,
   input wire n_rst,
   input wire serial_in,
   input wire data_read,
   output reg [7:0] rx_data,
   output reg data_ready,
   output reg overrun_error,
   output reg framing_error
   );

   reg 	       enable_timer;
   reg 	       shift_strobe;
   reg 	       packet_done;
   reg 	       start_bit_detected;
   reg 	       sbc_clear;
   reg 	       sbc_enable;
   reg 	       load_buffer;
   reg 	       stop_bit;
   reg [7:0]   packet_data;
   
               
   timer timer_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .enable_timer(enable_timer),
      .shift_strobe(shift_strobe),
      .packet_done(packet_done)
      );

   rcu rcu_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .start_bit_detected(start_bit_detected),
      .packet_done(packet_done),
      .framing_error(framing_error),
      .sbc_clear(sbc_clear),
      .sbc_enable(sbc_enable),
      .load_buffer(load_buffer),
      .enable_timer(enable_timer)
      );
   
   start_bit_det start_bit_det_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .serial_in(serial_in),
      .start_bit_detected(start_bit_detected)
      );

   stop_bit_chk stop_bit_chk_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .sbc_clear(sbc_clear),
      .sbc_enable(sbc_enable),
      .stop_bit(stop_bit),
      .framing_error(framing_error)
      );
   
   sr_9bit sr_9bit_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .shift_strobe(shift_strobe),
      .serial_in(serial_in),
      .packet_data(packet_data),
      .stop_bit(stop_bit)
      );

   rx_data_buff rx_data_buff_rcv
     (
      .clk(clk),
      .n_rst(n_rst),
      .load_buffer(load_buffer),
      .packet_data(packet_data),
      .data_read(data_read),
      .rx_data(rx_data),
      .data_ready(data_ready),
      .overrun_error(overrun_error)
      );
   
endmodule