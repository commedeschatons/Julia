// $Id: $
// File name:   tb_dispatch.sv
// Created:     4/27/2016
// Author:      Kenji Inoue
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: test bench for kenji's dispatcher
